library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package ApsVersion is

constant APS_HOST_VERSION : std_logic_vector(31 downto 0) := x"00000A14";

end package ApsVersion ;
