

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hIBbF+kq3oVaBXwt2/thZmZVCkqEUsrobKuL7n/Is+v4/IAZD+ZxnU18s3JR+GBgEFSO05ZDR/P/
xVqnh5V4xw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mFrbrNN2Iy2aMgLbmjyLagVGv1BRA/A/dAXtgEZvBXH1JsdW0tbqE7CcgD/B2t/bWf/vphzdyEfE
Qtz1a+CCHs4ZBStfoFAa0Kk2/N4AElHqndo2m2qkwB10dpRxHYBYIM8TsnGzjHv+Gc3MRRv5nDTU
c0fluXo+oor8ssR25QE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DijfY6YIFcLzBTBsFWeeH4jYfY8NXvmEK/hZQ9aT0hDSd3Je/Yj21LmilPHhv70y1trouG4tZlkQ
XpgM4Go6KW0FBpBt0/S2a5XkCoVlqKCnoc//o4WuX1mp91+H+1sSGdHdOtSMW4j5N7yi8fdf3Mma
iaJg/1V/iPoZ7fsaYSHM1whghXW3BgAg+uVNwDgKp0Xvr0+v0TXEnhMcvfJGCk7ZxZWk2u7a5iEO
OrSkH1tRBHn9Qs31Uoph/IE2TzjfOAWzb9vhqVCkYjlawx+iuHQsXxJdeZzjNlXERo16SR5o2JLI
GgcU9rsEUp+Hcxd2JjfSbszpWRHEU/3MaVNDkA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XNCwdX+l36YznBeQn7kiJlUVYGKrBB2zjt1UpGWFaIdIOQWhZL6zxzyLVbRsejTTuYPFOE64n48E
kMQtjnzPGZyr2W3R3SGB6KeHHUx9pNxyeNUyrOXfxd3APJdAnl9DigbPc/K+n0zkIbqWEydLVfIg
khTPlA/ncexRV1pXoq4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P4vVw8BLyUspYO28urZnMeeAl1C8jySXctEPFVvNqtg6Ihava9NSbOfscJ+47pmoPKhiyUWcqNJe
xZD0jdlH7PDpmGu9W5rxevvgidGt7SMfg0iUPqEmLLxZG6dlkSkZQKHeBdCxVW1l5LVS2iogdVV9
APcLIH1Hv8ySZWwT7HFfcdud0XUs4SZwhceaZ8TiRT3yp086kneb0uW/2QIlfzI1uwVMn4U5QPIP
rt59lNQNLmXYEhGyXeiqJ4sjMbP+3IG4yIeOFeDMhWUf6qgDysc+rBTvTouOsEPHvQarXNA7RtYJ
afWxcLBokJDKrgHjACFrQmNY1MmJtQUikTUFnA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 16080)
`protect data_block
PY/uOioAAACgRQiBo38AADpmM1iw3KPs1WjFQx2nYh3JBvmMnkCoCxSzoqn8s3VGmGeovhhFZuNb
t1TlDEZE4LBd9tfqSVFXoDGP37oMo0NPRqqKMxIkuC7WSucMiAgkeKecXMleQcchGqrfR39yVbus
YFZT+2klBK6Si6XcwSVme18MSJD/7mFOxPxEmou5g3tL4mbHtgJH1NDpWH8JV1RBG3a59zTLnx1s
iOtvz2CRUsHyTMkLjxeX8VSS+mrlD6LA3lj3dNqFCuiFzcljz3iz5B3Qg5Fe+q3XIzcVdtcO4sAs
uTHl/BAiYzjdzgc3eUFdaXnENbI63YEyJxe3TPqU2luURuZjdsgpJ5xsbSZx97lE1BlSOQCrwG0h
oF51ZgYPtilyo541Ax5IjK072a5Clf8nMQSAsPsBF8s8BJ1e0fA/7A6mCTAbeBY/9peq7YEko3HD
iQRKGuH8C991h/lLvbgO26m8oFTTDDy5MqKoZJdB/scEVPltivSf3UR36bEtnrmVDFlIYaOc24qh
xuhLSbBVhelBlLo4eBbhLbQBIZ01SZJMNs9vs4qQY4stlKOSm5JxGCryhjIduChr7OXPcDkcJWVw
3nSZ0GfDDCTkU1K/OvjIUdZ9p5/UoZNue40wfMkU9T1BcdYSn7Y2mCacAx7KbPCT+bOzp+Iwqfkt
PW3qJFFmkpPXJ4gZfA0vB20eNfm0xYNXT0INsgZ9hCiFoGzpTJBfpo4JqREF3kXa8wApaNDcaYOt
D9YAuBEwwQ8ntHAUnVTj69V038psF/iq61rt4GDXLG/cn040H3V0ERkkURu4X/x/ed4eaaBrCmHH
DeYNLtb0FT6EMk9mpuPVCxnY2pWNHu6iXTdRByuXjvzO3ME2/PzS522bqgpZfNNLx+CRtLB76U0H
keHBCL41/XazMg9Xhb5mcw1shMh0K6d8RY7FSYblguiUkrmU5/RcxYD9A/Cociu6511oeRge4GCK
7CgfmSAsG1QCElyCDDKtf/wnIit5HVx++PDMT0dJ8m5PXqRemcN+ytrezeMXncT9Xans/jHdsBSw
lBDh7FwpE1TlkkAPWIeBV6sRwNACC57ZHZtTHdAwa5GlV9aC50zo9GpeDv3qE5DEcXYKM9f63RAP
tHjpdJbyT/62EQVoPTLF8e0aq0Z9EZ67D3/AzSOfsIkoxnSzwZfxom1dBEkXeq89BT+JuYwsvUL6
PMV1f2qwDuziaubmcKkQU/uQXWtfgJj/lCnP3AU15yHy3VuaE23iobV1xf+EgxWKmLT68ayS+uGT
uqAR7H4PAdOF5EV3VcvQPOHy0EVvWg3kfLchs6CHOxINkkOnZ257B9iB14akW/UbohHAHcCukIuN
1et4DVqCVavUX9hAjwMbdRmMrHk4mocfpP73Rd87a1y8ecSvgYmiPVQmsA89Ht1BwSI9UsNfl1AC
RyiEKuXFMtRsipxXvwWasLmc0MJi7wDvtmcCcCWqMYKA1Y8kfqMqOA8q0gwUA8aHdvgcHhsFUeDe
pvDkknADlMOu29bwYuD3wSmAYWL2ay132iZkMzQfSb19M/+xtHTXf92TuKNG4uapbgZIEYga5/LP
7+g63PskO3NYqr2TruyaR6Cnb7ZYHUPWpNUNWIicFqdRcFNgZ8ImxaG22suMzf5f2t9m90jx/rXt
bVnQpiH0+k9apsbC/dmsIFMjKBcf0bIFbaknP1hpDDmMMMWsbpgGWK0eR8icIupXF1leowhfrXp6
Hy8tDQRCxHdqWcnnSnHc2oh7pFR8/t6ouKd8ZwomTyUG9BBKg5UAf/rVrRpHapR8I6quljq+8VH+
jchZBsnhbFO6FuhthxTcaY/PFBHXHiT0M22N2D6CiJOjEg1QsUAXGtl0DYzOIu+5c1h43gjESFse
xNDN2/YnRuZTlde0fIHdDlQsVB/iUIYencz82YI9pGJvwPB6FyfXyvgotbSuN8UOojTTwlK5hFkA
E2ih2ynqgQcFZaW/V6DddRYu0kM+z55bU4MZm4w01fM5ziPOqhzzu+U8OaCG5OfzhCPGsh17xKpc
qdBZblkiM3z/PGJeFXQqBRh3ejjDiYy+ifpytDyYtv63HU1q5a9W3R1k9KRT92QtUJquYWep7LfD
aGVtTaEp/d5GP8AixIVi1xmnUvGxgsK2O04Io7yMpQxilLFburzVMuMmegoBJ5PweyG4Wcix8xbN
Sg//+ucLtDJcb75DrEtnLDT4+JK4DT2ypBSomhmomUxTuEzqX2MnVLWLydvjTb2H9TbQBQdtI3lj
eKpbt9TvdhW+d0vjTW6xqrJSNQUJHF/34RZH+22Hh24inedfdCYrJ2xov9bjAZ5Okj/uRc4S8K2W
k6H7friiBaWlo+lDVlSzZRFxK9Kn0VFqnVyXhrkUPFAbfz7NO0T5HY79IRcTGHVjVKps3/MWg3Kg
3Y9Ats+R85okwmk1QACDXN9DVLMj2Gl+Ly/jS8fTQZrIJn8pqFWKlfK1uVvupI3dB307O9IaGRjI
/wxAglzLd0HUSoapJ0Vvj3zwV7suzaFFCj7Y9fkJOGVP0Tc0AxdRp4uDqM2+jGeLqzJ1X/9M45bT
wMKzLgnrHYNqW5FrPYkTssMSVuFsfmbMEz5PJHKm/VdviHese+zPeZknS2mcTPc5faM8piEbScnw
Hm6FbhWdDeaQ9X83obG/Se1/i4Ry+/d7VOlfIIYQGnT1fUly8RDhYkOnZoPXpdp8kzTS308Tz3/0
wsapfW75IRf0yYH+OComcVrbEuytkzuOSXmh+XHfkKt4fCRczyNQESCRjyUcHe26OJTIqHdpb42h
VApmnEhkDOcluQ3BfnozagFHHc/nxcolK8ZdFBzvvi5cF2pbHt8tRKBAjLX96+8V5QryLCRUZr0i
H2QQitZivhnvrFC+m5/C0CFVy9V0gtbIXMOSe2BhEzoOzZCoC56F4QfZ2i3i+yoEi42v5dDVWAAb
zPXXrq0DpU+h2kO6caEqqaRJWNpZa5Z+cBhDVA5/GeDtH6p7nwFiBEEanNoaZ6iGqsoZiPdXtugQ
bvC59hfRdwXwP0lmaJ/a8Nq3cNMzA609D/BK6j2Jy7EXtlidbCylDMh0PtXW4iD6s5dXHkqbRxwm
rzEHjPj+ZHO8yI4dvOpvUoJ1hYoevCyenSHAUQrMq5nFtpmQQZg0g/3EKIvtTXleDAuujufQxuNw
OhkP+SqrHLxQ6HwaIO8zDPNHfBTwPHx0yA14no7HcnwYFc9TZo5hxVtnlFIY/GnV4/A09PG2tHi5
ROQVHjMdnk7T7FGLKzwVZhwrBINUG4+Qwm+4r3rbNc2M8OE+a39lo++JYUXFaPV2EyEWxaCMmkpO
iBfcYQzMSLrbwF4G32GidMgMP+g3xo/YLbrOjIHx6pY4Kq5FwCqkmC8pmHgeY7OpuhRQDdXFx8KC
vkCI9ONba1nfRTtAZCtax9drT5YkXyKRl9tRTYRODG8h9cvNHrcjKWLenDzUP4eCmzYY8U9x/Ha4
ynC3/53905D727/OEaJhBwVWxDwWQnA5IeS5UHUcWWqRGMvkPI0En/XpArvS0GJ7sbOwsnh05yIy
V3qMBZq3pNjR0UFUoTycngR41m5Lx4kLZUg4fUiOUWEw1Ty8PCd/LxCmLHlJp45Iis3bUu0cTjRB
iptEempwkGAzHlsMJMlNtMahp96FVIwyY9VlpzfHMsxTw6TQCn+AQORhlm3G0HNHT35LF2KQcoto
bf3cb5KprcLed1aenCXpyy30f8pmrTqMKvH3gbd+1kfKmR/hkZQnV9ImQ2WTUifC4RKCH9b5YKZI
IvmUzDGHMW/r9vdJEUlovM9XJ8o2lRE1hK73G0UvTQzhDMDPpC0Xaf2yfDp4dfBXeSk4gHVy1HTh
8iGfm4iSPn72BkDl1xQ5d5VjDpSu4H12v0J44X5syZteXuXCrkiv56FFjjYj6hQlpUL+1IeukoBm
dKkIYg8oz+FojDigYEqKPFTQHg66BCxlrqbrY6eYMbz9vSntMJrw1mCIlkIBW8bgM/kQpQtUeL69
dnf+b5xCLFKnPcbOsNh/BwfPXbl2bjCWm4dFEIRCTZtEH0LWFPhVG8lgU/G6boP6s8Oes6q93cPK
DOIHLwTHDPuEurBhasBK/Dd+qtIpeIzUztJoHEwMfZG7dvc6WYXUfIRHckURs4nUpDuHPWa/U7pf
SJNM7Zkc0BoTpSl2E134TL6kUBYtFj3e8S+9NEqgsPgWlO98IxRt1hakYqnja+Fny02pwWpwQRBP
eqTfIJoL+8bvv3CCoPLNtsU09+qJPrsd12hbHVSqTpE+bKohFBwBBgi+y8muRyW0RdNeE81ielwG
+EjclBp4t8jO6w+Rc/CJzMoBmtlE8hCEo0zJUePWi5jyZp8mjyQdyXlhIx5QPQGVJgZXEGL0evNE
KCMMD13bvWMqet6AIRGoWGL2sbJ9vbDfmiwQ/JAfX9OfFG50X3O4Oc20sR8OxxIkFsqB4Z2SvwAt
A9jQJnCgU5O6iP89sZT2etTAleUYytE7tCwVVXxg72baS/7F0HMUEuacZT7up5rvHC8l9g77h+dK
K45aIdCqn9OcINcJD6ykjpQBXNAD4PbYvkV3RcGBYc/cVS6SU9mVrwMryOWnpai0sCToo50zvl72
mNbAASpF+WqbyI0OvpQdcbbsQYuLPLE+keFnzDycuhMXBea86OpgUW8jcdI6AKAzxVigwor0KJg6
ZnYJ666ti40Of3Ga0JPvDfvdLRHwGcRJUwGl7p+shZ/RZZ+IlnNIqNDl6ie8a4cEo7T7ogoCuw82
fa9gTH3zsTaADitskUxd0qCowMyDrxJWZV81vO5wVHQr6IYAvR3epDH/EtPKMtrEbi1pp/kgJwhK
Q5odUvTty6MIsaO6U8nGn8CyIzYjzd0QP0djeO9EsHg29jH16rvjsgKlXkQD/NHoxWWjyXoVfpCj
CHTGgBLizIYk+rd5QG3Ob0lDKaBrxv5cuswebdz9bg7q++G1xrUrYVGesE2CeGEvGM0y5GztpBVR
4EqpxLekPPsce3pR50CxFOG07yWwe8BJjXWL3lbEsqSwqaK6BoXCbreCugVwrusjL9bHFwqtv5ml
h2IBh1BkbD5ftQyRr2y89uLuxe2/+18849KFzPPkSA2KNuqVK9e2Esl3jb85b4qzFL3qjEWG5waT
ZO2ufRAUxZZ+HbS/oUeHnj/yVlQ3Zl2VS5VroLTbcIniCJFp1olzeqAlYGKH9G0ZU2ooHjW3J41O
7JoRZ3uLQ6I/oP72LEzG/RLW5yK3tPUvp9llHdRcO8/QAnGy7Pyvv1bQI9I/mrwnzHK3aKB2QZcW
XUs1SDtt8gkUNBWZZHcjq2SH12UqosCSjhZ2wKSwveGWvL0MO/f/4sdd8U1lYN0f5OFdn3R00YPw
qkPWCxdl8CBiNdkA9drZVoZHHEyyaw8zY8fJNvDI0K4wAXBR2MKmdgFSlBYbPffuvlvCBPggoYHe
wlvTtR7apaUFU4mqeeKhzQizy9ZqKcuMyvxvL9k2NryQJkdTb3jQztsi3ggqUIJxt/VlnGlM/RPc
jpYm7+7/TkdPnOxY0fc2GhdFwAP/xFNul0iBXO3GuHtlXN9/e0s4VC+/C1PUKgPbK4rhKMQadY77
berd/M6WKZpyU4d34Ttj5Bj/AF61bCiDtPnGnC4QGuSSV3y46aFlV9EQt2pgzU/J8GTvl9mD7nmQ
/qPWmdUdb7SCwYekEW1eGgO/ccFaJyMeTjAvGAEkxRlwWQp++55D5BuSfCU/Rao2v7KkqUzsiWLk
Vs9VcaZfZ7NzArJLcvMgFXG7x/OwtlvDRdTlQE5PKWz8AJb3/64A/n4Z3F9ivOOy2U7TbQLgxjAv
8LET+Ewix6ii+H1K6PhrseVxI2BJv2cbh/MDM3Wc7wi6Zlu12d9QBSfDuIgkpcjeuvR/E1FNttgS
iZ9AmfElKqoiQW/s9HSN9lZSGXCwcW8q5tLdVEzk2BDuVQPOEXTxQNS+jYPH+8DrxuKvrnsfbzLf
7CgQ3+b6mcdZ3xVXg5psc6Bgr4SLv5ybhZi+kW2bewmFSdCOhMkf9AG/aKwQPtz1FUaOaNj1B2tn
epevOA43QMXbpQQWNFM7bx+0lexHrlRs+uWiuNBff2vU+EiYbJMCHCJK9WsyJFA3ncc4tTxlVzDt
eXrjlrmk2+bfqXV8CVAssyzeWYcCMc8jZUGvJCOk6vF+8GzyYXFDMeITGcYCrrpaX3IC7fQRE24T
/ta19LHQnQVZccIPgdRSqoo3n6OvCqDYTi/FsEQ4nj1f5+SR7wF6JggFJ/S0QrlaoW2AG1fUFju9
Ofpub6Y7+O9+kpuMlRIjTGdPFl1rBsWMRF6r0JlQlPpoTy+S+XgbEZGZnH1pFE3f8h4qll7p4+vs
NQChmNlpIvtba/ZwjFdtqg7VJiF/2NG2vbE6i/JKEm0aIXlM95P28MkWseDoe7++Cguc3g4AXkal
i4o9tpUgmlnQcEOTHhJItxdMaIXokMBq0HvPUWDxnFmuJ5tTulAC9rvYmmDEbuQYP7oWfFJ4IXIc
529fSP5XvCvjXrPqpOIZACQ2OBnZfd3DlLpvxw1obpOtKkxyHz+jKzRgULMStUP564qWtWI6QHLT
5BzdUf+OWCyKoRkTdth6jYlymN/BTfmaeRxluyVZGedm5yXZqSa57eucvzEE8NpS147zmqxVzJ54
QAXnZsonBRIIn+xaNakHMzhtjcpbhmgmeQC+xXOqAENNEv5P8wSMT/NLLtwmBuiuQ5OwiiTZtQ9L
lPyXpVu/1Br0nhdApxsWQ9kKVX5Aje5AA1GDcJUHU1WHV1pdMtcl+WKgrThIJEkGXBtcYlYK0/uY
ksQi9o63Wu08mTiORPy4c2iRsa3edDO/z38Eq8CZiWWcvjIRcvFP32aapYjGcuFYonZn0xiMSSZk
7SHckr+QRiN2UHLmvbi9xmP5VlGGpb3AhtmPUg1ro8Ucr6tlwpYX2kNIzA52ECxOE5n02ATNU4Mi
IhV1kjw7f07/awzPOJGoXPkXHN/vAkn1fUqvKBCXaJnZCGFidvfyUmDuRyFnoQLsUXj7Ee/AMxyP
8wZL4uWkyAl38zIvWfnfx7IrAm42uwiTGT1KjKWUR3PYln0Ove+CTmslIr+sflPlpPGwuQ0JaBfU
aAfA6y14Ywcv8kY2QbMv1PMh+pRa8a73QjeC+CZCgJzmDYO/Ae4brJz59OnyMQdQ8erLVbzYG1pz
omvsoAHA+0y4FUj47ezGInSjxgwgYJ9SMQmgvDUSCWyBOh9o3pfER+LApL1tLhe9HoMByfyaUgrW
IgJxm2vYre+4c/BIEx61GsAL1G9WHyfLBi4eymBHVN/+5zZN0Rv/1HwBnNqDHBJQQRVOpJLRgDv6
ln6HcM3nhP6J5lhbWmG8B6fJltma8r8IGmaSISu5SMicz9dLc7+mKktaTr7g6qmm8bdq+LrDXTVb
UMMyLe0iZnMkDxRrEJaaNJOQ5KRwTxG4I+cA1Pk7uwOeFk69Ga/359HzQzkDNeI2kFh++dVCACJR
k3bSsitaeZqMZHbz2RNrczTpjt0KGhIKXtlYLTQtu50V48p5x9dUbNk8Sq6WKoWcpy9DBOXgDjbI
d6+D0A5qb6HoOtwHQmM/YyqtyftBL04DMamHAhXPDD2KV1VRFmaoF0OMNGRwnEs1YkLSLZ6lXkm9
bPDmZD9xaA6iuXGS4dk4lSfYb6fO1jswa/i1C4PWkaeIUsSzr/kY+74w72oDz62NUmvwl+lCXGct
ynVM7SYpt1HGBcfNWPfyJTIZmOzvrvJjHle07sYXFEDtybaYP8c4qobmoH2WS3QsbzovCPbSk6AT
J9jFA73HPoBqlI6q0C3Il/pPVcW3gHdt8vfo9mBRTQr0Lfqk6XhRhfO8Yb6zW+VfSMZY/zy+SMtA
T9TnG5DPdpx767LTvGuc9eU7pgXyQ176swhz2inIK/Qq4qiLDs/E6tHIkmQUoWEXp+tneJD6dWqo
gwk3A7NGtK03DliymOhoepfR8fLba/cHsMgLW+KeepasRTtsJkTqRgEEkeSFlT2BiPJq9vF5/9wL
+uE/iGwvxF6KI6vqqeAj+SUTCLsTZ/YsQSWOB5i6t7OKQyokmMiYZxV5miZtzOhpYokeZTAJIry/
i4l/+u1zfrGE2ysv93SIAia4XlqE7ULNqJIAI0ahwSPnJLDsCBOha5Z2lCtqGQ66sDgmi+4c2pVU
lfPc8aq5O71naJ4YgLqBhUeCh7735MABxDaR7b+sUo60n/bEWAm0DbazRJA6Ayvpao+C+M88LtWI
hrl362xO6+yv6B/LaQql3BC0xfgbM9dYSvIklak2KL9QdOJ4BRNLWQBB3hZ9ye03TxCoGcz0YaYv
VKY51rwuD364wNJ4BHDo6Pyay9GKYWQ35zJUHCSAGpp+V5D7A5uCa4Ud2Hh7Kq7vcW3vPorFxTfu
2fGIpKyoE3gURzhBGNBmW76YS/kxVvfUinqgj3oBqp1HlHgjW5pbBOJ9dkfB9FJacZmogW+gYTcM
jzA4wtnbnmfHVOYsRHSzwQuoKByhWvX4t48Icz/qR4RBUHxng015HMuH2hFoT8V28SlNkkr8KuDu
UNiPbN8bp0/DXV+IlOGCkl8I/361zQQ5f/VvM0rUZcX0MX71aZyLiltuxsIpwGW+TbbK/sL5NvXa
yfL8aXWOxANzbHVEvVVfA584xGn5WAEVEDGsP2L7iOOiockRGn9NTQksykqBLAW+OmIVXHOd3xAO
HtvDzA1sN+ShfsQpqEaM1PQhhfEFpJAv8vj6NkpUn5tDlH2SLaRAGxfI2hTrxZ4TMEtftWCyIaRh
dVS5+68Kqbgc9p2p0M42mWGKZVgsBx9Pbf1qd5V30BoDp8CgNHHurP6ZjImIFdcx//JOS3S6QPhq
xWnhQ7VnSKujUeuKpzLKaOvF66kHLJPfBybLD5XiZB/Vv3JOvgeRsB07yKwTgM/4vm59QiytDggI
/DykdNimN3Xyvqa+vfVGKPfdILBm6lUpHweHYogBDG/9drtyBPk0wgAmWYBVZOncplTh2MloOV9N
35ts9bbQry4aFW4lpM8cVzdu8GF1hKkbxCimvf16gTd3BX1eS0DmuGL2IqUzoU4YqR137hBCG7hF
Lba3L9eSm/WxFvE8fvqatA8YM//LiPU5Xzjvzt4fVbn7YtQZnCaAV1uIbBcuxPjlYvWBl2Pmkt0S
hsoZ7ro2wI+xG1uEPcfoLMzWASUNMA1zA4KsVMHWw+raP5BoW89hMSFrjo+daY8GqRl/P4upSIhn
CbSddXgBbBwkFJ8jJSOnIHB5Ll+/1t2NXEHRjgz1gUae5YjCIxELTjcQ2D9hNBgfe/52l89UsNBE
oNR4gWsu9l/UmpWSOKjpKnGvAHPvHIauF3vszxImFiOT4mP/p7aHnzPbg88tpl7zomMiEb1MrWvI
uJ1K6t3AV+cezuWAMH948KLXNGTBM2n6XTb/KoiMM4X6/t4CPbQEtcVhCZy11WWyz+ycL5uxCCuY
ddD6k0lSDYDBLQ3tlgmA/YhOEZoqVpoFPm+5s7wzI34bPIKRzOxNd1Ug0AvMX5QunsLDqSmMGqY/
vOQYi0ra45Y4hR5yKfVuAklBHKHaXZPyLfaT9cYZnk09dOJNiM6xH93xypCKiAGhG6TPH4/EgiC+
l0RtS9eZdiRnBy3f73nflQBnsbcGessJ85DnzPq2w0WAxdll46tNlCTt8B7eRDvX92BOsVpuMxu5
654Ag89vd9Ek1yaPXPXyCmnOQgs6lHyHxWcyYVUfQUVDx6z1+Hya7jjvPCZXnEg4+smzkq8Al2Dk
4zMyvmppt04GemENPUOv7ueF/VfPE0ZAFl9FBQl9QrDVRrglS+c3ZHIAVnuef3e4FrZAx3LFpa1h
epkEo/18oGC5LS5sIxZqpMqDv3TGMk36VemNBrVHdsrr3nQyDxAbl7e66g8hlRzabZYyk1KHnIym
fS0WnRdslnPM7CJwylxb2Hk/K+xmfW03keVx8m0qY9vwvZG4jIwyw8adIonXBDG46OLJUyBfLiv4
HlNdbsBmWJAP9EIrtyoIOX5/y66NjmddHRoFiDUIqGYTVlzZRCOcXpX127OKYvtgkODDVxFR4n6w
Ah6TrsljwqGMXOZoioAiXttcjeZmmr9ZhvQue1CcsBHC1AuMpt33VMH1OnOJVDcpNvHdaZhNrMfl
WgdJwuU4ub9S3qNQyNiguS40EDKltVqzPu9K5GZN8PY4mE7wRbQlQfVNvYkMOlXzGAFoXZ0Ca8kG
ryaYJ9lZ0V3ykLeV2SbH04RhC3TTerXXbqfkXkeawtMvq8NT13wuVZ9KSnPcj67lxTCEqnhdpS8X
GAW1c+YoUKBZa19HPxIRATQQr0SsKVZBfhB38UwMNaCr5iWO0Ln8YtDvQ4XhMOivcAwDh1n8S2L/
1fDBp95tz83FuICmaUg697QCQjLCjRQa2WeGQykiblc1Hft+cKlWn77PHiiwGsB4HY3iPLImkVzl
VWqr/Ngqz9VUVPStZF5FmtsqtOEESnZVN0hAox9G7Ej2ox6V/onV2w8rjTf018azU/zGtw6jRHGy
E2PrqNxLaaBo3J3rY7NcA+PlTsXlsLreZj2rQUys2djG6XqTNxnn8M0IhDCg8pWlZ67GWCoI1FBC
xaVyIMIw5i2kwXOh/hzStRbJn4c/CZc4gADmN/ehk0yJvZ/2yKUyCulZj0sJ6YmvamopwjpWi0RP
3KdwI86kSDpYbQm2NMGK7N26cYIlmPO9xlflAJBTuDvCP+CY3lx5d6vnkpYWh7qLOpsUVN3lHtiM
kEc0p5TzzeolM0+3Njp7G7tHFAsGoMY/Tp/ll8xPpBY+GCFBaNmR0cHh3niM/ktHRAsr/T/9crtN
QGys55aQcFwHohte2CiYj0l7HbxOrNtHWDTDL1RrQVL2IHOh7O8I8BMmwc+2tRqUNSkWp+67c11j
XT2pBdRsQPDURgMKGhqlSJfwpseqmUnRgnbrMVMJHOALbwD49TofTcCgxL02Avisz5EQo/UVUoDE
mzHKA278GZ/fVDqAO8LkV68cVLHNV5dovBx1zbn6PnMYPIKp/ueLm3ez90fHCTcya0027Toj9sW1
dymFha6h9DEWh438uPyoq8rr/3c8JSaVhg7YqWA3h1Yjqv1g1cOo8Kb5BTD7QvehzpFJ6Hs/u6Vd
EvOYr5S7cJTLghGGck3XiCFOL6sGRV48m/XebqAWYKhRnkrObaR2DySz6+IEm8k7rY9IC2uWdDty
taLjTvbV3aFKnCE6coi2L5seFKjcR4ihx28bU7VQkXs6sOyS1eMERO9DQ1p1M9q4+ol3MePhyPUs
pXxOvO6fMsM3DnOMHSDyhfV0/lrq0nti6PFKt7lBXOhRMPWyr1LmMXrtMwhV0cXA/iFBpIGLdFcF
UTQuB8NKlL0siyj6c7xp1p3xk3bDR1xuxg9Bg2vesTZUzXAEFLeSmQhQ1tw//w6OzuPd+B7BOAtE
GYZw3NXGL97f9XhQQ6pbwY8qhkCrE4f4Sw0GFm+ekCzpSA3n5iWS8Jmg2r3RsobCZwquu8lNejv+
7iexhMV9dIVow/vqfoMkgI254jG9FfODgSdSjxZzasienj2XsZ+iePg3ad/fQU6rpTVfAZouSekR
mrPNxb0iHhY2IaH6RyPXey2shptWWkBbNGhpjB6Muz7xp6KG9RKoBOheDsmXfaGwqQKRwv5qRSfD
NCIT7RoG9WKaJsKK8PeGbKlzmkBYbuVkFyVFkuS4z+4VA74X7CwVhtioXTZFOtSBmve7ffGYMb4C
p3+amOZRZwa0Yo7/7k6N4o70QMlzBWO2BcS4xSTkHpRfPh/vZbfQzUBSYr4Yd46Z7iQUiKUafN9a
GhWyhFbGlLah5uVw8e06XdEEko4LmW/4NJXsgX+1aJ9ZbWfJWDEC3Jmwy7Lvm9v4juaKqRze1w+n
DkpCHsh2LXA9r6ix2IAZOjF+W1XVXz72pnoq6nxiMQ5VWJlDrGgGmZTnG9x+SjwUcx6byycch50f
HrPJ4c3I7iQHgGf94S6WYqBIep6Ot3GYUoySun4iV89qwbyD2kqf3QiT+p76MlOxD11IvZGdQj1O
/AZfWDJKmPDWIg9JHcmwh0qbZiZ2Jj721wThneHMhCnaVmjWFBrh1m/0LkBBKPVchWYrbZC1Gdoi
CphJ9S4m2lddpyQvmXDl2kY/jfyE81fNmm5yYQz3A6iDv2ZD/0e+e8yBrgHURxhPW4gXkjA5FNtg
4kL5hsKoSObI0xrqWsM6bSVc0ohJfX+RQEwDN6uCtL8FtaHBCX0lpaWxNlwd4x6rHq2662N/7GkZ
bMHnUz4EMjz/kjYAIJ423BW1NrPCjACB2VaPZEwLLat8CMJvzatqlGJ2BAZCRo4iV3KrtWte/Kir
L9FFFhr5xNmaS45Slpr0HopYC/+JW9C4FkRn/JUoiFfE8U7f+9S9tYFMX2LufYMvz79B7mXDxsrG
IKRpki5UADwq+wBrTCRNS0MjjIRu1gu3LU66QH6gKCLBg2eHU4dnMo3Ew61NqAGNm2YKk6dVw1eg
Ji2CxnJF2PbKU22bG3f9kiensDuZXT3u4AQHn7GtQ77JzDUL36ruDGNQpa6yQNZ0/8I+czd9NbPw
npKoQ2qm6CwXqKQ7VPYLsFwgo0w8VOq/1C/st40G9z5LmkAMMhl8kXeOOGIjYNst+ATin0h2Tuul
Sw293FTtcYJzupAG5nRpIhiEGhZ1SSqXoE4npcS18OjuSZ9hFdTS9eje++k2h4nd2vchHwmzJeWO
BFUAPhDAQv+f520JpaSr3HiIZCt1JV5q+vYviNVFNfyQmI82IUclzpZ+sZfL8V8YJdE0j4XMNuI0
hHT0EOXbec5qvEih6WSWhvfeJQA0aAcUHit6S6OY9i6ZAm7qd/bEjpRtpe1GE73haNaxORBhkRRO
lRqU6X1XZYCumAVrubGpGrRFEfjo9Qylurd0mry/y9lCoHK4xaqRIrzLhkuRAlC6UPlZpZCEN2TN
J5c9p7AvJ0Xrb954wRUOfwMT6Gd0bUosDhzM+2ZQqQd8FP5hCyJ8vFt9eqkA5tWSpNI+PPG1vtQz
MRaTB7rz06tl+Tfc0who+rqZABBfBgUk2fLntasB3/D91g72xUd1b/zQsiZFf+RfEedVNbQ9s2iG
uAGT5trdyfOJoQfWmvcBXcJ2VqK5aePQu2Lobzg37FWwp0sxr/XSzoVm/t48L4rRgCSTAkzajn5s
gY+crditoukknooSwM/8KngqelZGJ/pCZqvqN+z6rxp24FgCl1nVYdIBxSxZgF+/ovyxZ/XUe4B6
MVJAyZZFLIWQ7UVGkUJCIjTsx6jgA824VkjH13cq5rHU4I9wn/MZZw/gIQAmAuRmB+el9MBF9J6v
9zxXDhRVemH8PjQP2/btMyj5TFL1Pwht4btEOMLWav1VUfP02AQ84uvxzttGJTz41htF0dT5yBjU
DLoXc3bGjuiJGJ/jcz65MT88+b6cFHWOU/05iwEufGwwQkQiSnnLLVmxJV2rdI5MV58bVTIupWSy
5+386qqhOZimtlbQ+P+2sFJIqrvm8y2459shxxo0Ve4MUY05/x7QQ16J7FnbLCpm+tp/mn/aldVF
Ek0REClYHbrF4RsB1zedD57Oc98c9Hv3aVkqgk4D7WzzfiuQKS1krfSUzVVl5yHRxu8xdqgKNGG2
PLOT/S99OM3UzaJRA/ia0WqeET+/oLc1RDYOCg1wgbABRi0Pv5MqhNovjBSwDTq0Cr+HOH9s4THd
D1QT7zB1xTn5u/vBn9qkBXtgp7LlID5+Jpin1z+CIhr+ML7bCgij8tvZbgPOpl0IB4pem/CBVVkr
mwH/MSPQowrmvQ1EgzD+5lDTNdlbbKEkl57q5IZUKzUU7rP6Ju6lv0zFngcVM/MRp+Peq4K0k4bA
IyZujDLB3hs1cmQ92la5GVucrU2FE48ARs8in3lWQLQ23nN/PmhtuATIDvpnWMIzO9vvq57WU+cB
GcrbwQ+R0TedgBDsTq+z8CVzHSDWybA+mcm9aXtjfQjsLSmJQ8TXs5MVdJ+S1a2KrpA0vd6zD7CP
jtbNUqLNqPA5KBEuJHV8ImOx0pEZYrrbm0ZYWxBV8Nih4ZYJEPZPWaPhCE3baKYIL/br9cD+7DD3
hy0dijY/U8LNtdJVawy+v6nP/4+PpsQ959kYFy9XDQ70alUi5jThbTy6CL8kCsvtobLnMaYekgE4
9WQ/pcNE81Ogdvt83jHyMCtUz/1aqFIA6FJZBZJeGd7Ft0eKiIoDGwkNkFVrz4rQn8+xaXS4N74v
lvS58sk9HSHLsx1W+U5osx9c6HqWoUOdXSq+EFYdbIrfXjGiSPduoib6uz3puWdwPnqTfMZ6KC3T
1sWQwnhf0Q/AKx7igE3/ya0u0/kUyFAQ5PaXXvukdsi+kj6uLpyrSiCpooeGaYiVUzBQL8fyoMhs
R2xGCIUfmCfuI3TiPWVSMLwtQ0zk9p1okmoTv7ZxklLNwPYJI1rzItwBvtCzwBkzkM7vs+QOpZUP
GuX74HYd1gE5RIcEAisjF7IBlZ3t2SvzMMZf5tgeDp+ZUO3zeghXa2Q/RMi06h5jklpWyF9ItZaD
6Zfg4Azklk3vR5HPRF9eooLKgdjmnEN3Pu0k7VXCPunGzJG+Yr8KYgW1wXdn2xFYFFro8c8aUL1l
e6RhiFYdIFCZ4s6blsnCLIZbDpX5YKnCgYPgbXJJwzGZWt4UahVQUEXWnhW5XIXd9Gjm968bpC2q
L3Odszo3VQjADvwSYfmg4sNyR/UW5/pqqDaRXOfuO+UlRGqNcNNt9nMjFXhbuREVPL0u2Q65VIOs
AiCBbwDIEyRqztaUwCKWDxitz+ODfSqdZ0njsoZN8Gvc5NIvDbBo/moZ33cQ4m4ojE3Kr+hEBntV
XGJXs6bIO+uqAAaUW6yTWswP6RR+cHziiV5+R3wa24HjjHj3Oyv77QWK0e7yoUP0EA2Z3fNlLMwZ
6enWAXJEOQdNgGUE3xoC6LY+XW+POfOFXfP4qM9phcbyACrQ2MkQK6GLDmgnS8pvS8ipvtJhOspc
vRPQXF/PDLpmjzSXsuDVyZQH5AXZqpyPCn/BjJpbhFjm5+cLXKWovdy9mIo/LoujVekzJhn1i6tU
UeKD7L6J4D9dlFc7y6fFNIT7UhLaXBXZvMZNvahFGQWh9few3/kl2+taadcg/RQ7ySFofQXmxSHV
NGINxsxRxLS78kMuTEM4Pn6HAQwRoehF/eZx3BEIlfUseLh5KGW1v8L9P2YbC/tKTZtjWdQnMkpz
dpL24SgvIX9S/hBeVIe2pR0NhPauotiDcDNR4oUZp5nwZNXWaSnwknwn3pU3dT09/87mSndwxoto
9qZPsn9sfIJtod1FnLWvXGUbR1/vWMxwjUXDwgahIsBS6G8FxNJ15PH2wklkzfZtPogHPBkCr5BT
THdtXceXy4h186YPoljB87Ux5vBpgdPfUY1Tvxq6suI8yU4R30uL7qq2sGJ8cGZaal4h+WxBravv
nigQs/Sd2L6TgMvFxNdp1WkWhpLEdB+f+QLpliuwefNg8fJBkov46KUaXtwjmmO1BMqssvUFzrBV
fLVM+yK/ARR1+2v0nrAUFzisqSRDog/pf2LjoMtkvhzwqcS+gabcp1CL/69k8TWCIl/3JIHKTBw8
srWsE4czo1bqJFo+3BZDUd2T+e/kAR9MgI4KlnJEKxRQO4y0fX/1sbp9A8QrgWTMnIwL6FJxfqdl
Xcv84IAkkyakKYjAa1Sp+28ftbM6LSf18crX9c/W8zKmR9qrcbG40U1DcUgAEpPEyGrAC91FvIoz
yvdtOgr11BA4r0Qm/FU8QVMLrgYTJ8XeuU1ve/HFsMKveupuyvDrkUd0vphYJXMQx2SvTvd3O4f3
dYM251L8wWYlQi/uWBA1s9oKfvB5UyIm9WpIFGPT1/8QGDpTw/3+uUcEL56nrSbLxCtuC/EcJ8lk
24foxwnetJtzuIA9drfzFyM2a3AJ7uMsOkdcu1S5iaZRkRxeDqxF/a9ObkM5gxfhFBhTeTEBo36Y
KxQic47DvP6j1N3fL5WCG63mIGevZ9TDW2xme4bOxWenlfejyjQ8L5hH+mB/A74mtlK4Y2QRRunN
3OC+9z4MA3FC/Jo/RUpjVI0hJHJ8oPZPGLqn1v7we2Q9Ye7Y+6/R3aV3Ji0EC6tbG+z631A8B8/j
g3UpCTlm05PbImdZUv8nnElV4yTcxRla1DXp4XBsGuJ6/0EXKbHTfbKB6oioBYMBhjzUw6i9uO8L
2Dpap5L3YQyH7BJ/8avQFtkDqktwH7DiHBCRLd5UQXPMQc43AwFaJ+W+c4DTKz+KuArgdLU3E08U
vo06ufxfmoR9fy0T/r/TFdnmaxv+pmPomWjlU4dU05vWGZbmZMpO3okYW+lFaLCIl88qLlbMseFK
eeoSvlFn67mPy4cGX+MdxhqHNBycvItzhgywdqAuNuG96zPJ5JGrvnWRe+DlzS34QCvF2x647MvU
OWSB9IyfXmy6bJYHYmaoZRyUdQsnqBTh9cl5shTDCK2SEXeZg/PDzFVtmiatXW1FgXtQE4LviHpi
jwwifARRjrc4A3V2ywA4qsRKGliLGE7iC7X2koZR3cdtdPRkiy7c6XffXHK56UFNF+hrfxlv/5ey
pJqKj7v3OtHd6vsrrDBJ2foye0aVJm0QhsmEI72fDIYLa4WEhm/A9ND+G6dmnVbsPpSwuouniMhE
BePZ7a7wf2T3DYVj4+g8Zs33uj71IDP+TdIGz2UlQ65DJSn2z2QOlsjYnhQb7zbs1PiAleQyAMxW
XyxPwJIHaCRVPNlUEvWfcK25oHuIhNioql7vuejvr9GhSOnoYHbpJuFZL6+fQ2HKNXEXg9uHI+m3
AB6P+leH9EwlT0QB9sO567fzY5t7Phf2xOb1AqCfeg7MpXkzLKTv49Yp4PhgEELx9/bYiA3UVKwQ
7OipTygc/+IhVz+NK4TB8qIgfwglruPvQXh3FFH8B4vqS9ar9gQQ18nL2FEjuruzwTIeUzUZ8tKu
pX1rKJGfcDduFcW1eK/yCeDnLSWcWlUFzMIJhyv5DLqJTJfS0dPFEGECKoJLB0eUuU0rBwEDlUD+
fzPlOArt7xwRa2JljPlBU5EjK2rJv9LUCJ1iTV6clME1Vl/X50a1dgaDcsZFZg4ILQzE0u8LeCkq
hJcRLVeWWG3qCBI9J+dfrMxzSgK6noT3ccu1nQQ85xAgY0p6EC8PxnxnM8Vf+6N1xi6R8rCCk8Ve
yHeXMNk9m4gEThOB83GpW3MNuOkgyKVNrfxu6Ix/RcIyth+YGycTa1gr76t1uu/XgPJJ/OwuvL3d
y+VSLFWredvrSOP/lxUe4g/2Ku5g/0Et2lp0/oMkzSubjsWtTYdHzj1GS0hpFjokI8NXWe6tpPEd
hEi2yQ/Ute9fwadoeLPorF5mTAouRczkkr5WylLUpf5dZKiTWrMVRv8qZGuTp0FamckNo5QJ10v0
VB+tGyJbBfWJTb5jzZX3qkoitKE1e0KnV4SAtf+SiMQ+PtL4NmnSbJmhVP2oATlLZaySGBf7g3Qk
jdZghsajyEU4cvVnKgYL39Ko/f38ee5J/9MfOFdTMHLekJQbtu2NVnLkTiXq1OhrAAs3ANvuaIQv
EqQAfj7ofhjRnWbr1uyuqNTVfpnAWBJKukHkP2jJQiirmB0Y2l8uG7zeXTaL3yumDW4WieIXxJXi
kPVTy2m/jn2K437KIpOzWldgZbaXw/B/VbEunb4HTB0VhYwuH9kJIT/Y8mpVYmxW7jqqionJx/aa
JJ+WrYXK0AZZXRPK/5wGQXJbppXJ/mGVma2UrAyGyp8tb/K2ncK6X39AcesgzZJeQp7FBYbjFE1C
XOyNKPsHwezp870Cqc6bJZruceYm3Qxp7ACqqn7R1+gd8ku2KFG5rAGCV+1OYIQjPa/Tj0dSmYYw
BEQQ+OcrbcIy1x55CbW35gPRrG3tcnqH80sTUVR4dJEjtEySzpFJxwET/CYRZXjEdv2pH+1nsZ3D
WAHvckAhmkF/OJFPv/d9PWS2wdepze3bzxgYZtxR6HDSRahBNkz/mN1wIcNgxVMysVJcGmgpRweS
n5oewuqrbGgw9V2qTSCAHhdQXYOd44F7oHdBFhDYcGaF3iNaXkCRfp2qP2jZ8DHCTDbvMKgK/hHH
pmtseX9E1ZkWqBowMiIpBvWHsWQ6lZOZdPulIHX8USNR6xPCeStWdSGBke+tp2I5ltb4/0X0nu2k
CF+4YgszeRsMPAx7w1WuzMwblJdJxgo/LvK6/wMrm/FRN1VGQyVan8klEZyYyFm0FWPZP1OSdNxj
RFjVrdCWiJCLf8o02yAsRYN43WD3YRRKKBELKdCGViX6HZLhx1+rUYGBnXeSU9fhx2LsUI6IN2qu
isQPJ1C1gX+cKK2Imcrv5TV8kcef0zJEPzwMpYWhSiq0uDFmWMTX3nXipJSZZqHrHhec4bamQGag
G6e2vN6NVMJxVw3U5G5F6P8nwHycKfylztzD79ciKdRRnV75cooQnSrN9kFWL3iioBT/Lt/zjnyd
6XHOzoGoyCcN6Uf+3HIS8SOzbTkq0dejUwbwVXmEugiMIFQ+TURqy5B3QA1Q1+mJjgv2NEKRAXr6
LZ0CuI28F6DbdDMnRshfzqegaT5/nLYnGNPFjYweCOI4OLCMjhhY+fLEil3ZtOwP9buLHEGChMj9
7kQDx7hwHixtQ5stWaRhs/kNgtii9GzKzeTqw3j0z7CpAzJtJXWwrX8BmjAwgsZ75EGqB2usIlYs
QI7OQEkLLXwp/Fi6IVARjCTGP3oe8CUpE8PeEGIVg0Zfw+ZrFQLpg54t8OdF4bblqkVOXU4N8ovY
b35U7ydYSIeZkKudBXyu6F1aDYr6N/6zgaqnHjZ0fRIQJoPYYivtFnHDHX8TfK5nTaJfnbK1QSpt
+i3dW3ft3DB4P7s2jGxNiFEFFoigoc09ORPIdxnBJfAa3VJrDGdS3ITVMFtt1ilpeCaB+Qhb9JzR
30dqVqxosp1kxCy823AGZSNjSGMOkWydYpz3YJ8/UltFfEl0cbQLMjKDdSt+HCkFZHy4cGFJKXBp
gP+Mr06c4DLiSokG9P0C2mRNZWgqqcNnfVbbn7plOwCN+M/PIKRRzkzE5l0eteO563DQk3OtR4zX
6ET6Hhxo72BAQ36/UAutjrzHCj8nUvVldZd405v4+ZNKMCmcad9RmLudR4UttcuKvX9Q9LBOatA4
RGaAaKok0TXgGZjyjnRwXrziJkQrqvi1WJAttaRFfaE+NNNrueb6XelHq3WXlp+2OVTpuaNc2NJP
7caSbA1TlIdnIG4nLts3FSE5o/gOFOmDr847tWHmatFo7javEd1eBn1QV9Yf1mcGF4cXESYH6qvf
qhpfhRNW98k8j4VgxJtlNrVtVdLEqUr9UiB2WN7wd102z3Yi8pByo5YgODbN/Vq80ZiPsV992oi9
NilqCRBfVc4FLWXgKB39MkfUs5QDm4gdIUih+7WVEEyt5WWRaK3MKI5rW9gyxmoF4murQbM7fEX0
wfNpxfy4PXTj5SMMn4TLWigl6B+viwTPt4fVfJl9kxk/lFSlDsEZedfcqg5dbwsddgswuzGn6Io+
QNXo/jJTtaCr3SaW/UMHmUReVpKL5fjL5wur2eHZtZUmxiRzRJbEx3K7lv7G8DKJI3PPN6LXNe0p
/619/yBt/NHdH7VjSxN9nzvcjwM9a/tVURW3mTWoGeCkRxBDCP2EVukZuh5AJBLE6OVKMjFGK+E3
srZdqcuMnUDNEhxqwdyvOC+ROhmXEPjHGNZFmANH0paYTpU4CocZV6M3BD2KC0PuzgXjUWkYyb8Z
jMutRVyeI6RJ3WpdfuNSn93vaDaAvdCDQ3T7Q8FtlXWDuybDI4BPTh8hD/wtWQ+gOwupBqX8UCAU
gs2Wd6cNL9ydTJq2sJ8biAiW4VHKC/1EVQtCHRiCniYVuqzrm6QswurEEP3L5HlRSLJj4s8bm9UH
z9SZD8QtyLbjIZeLaXFZxEdG8AMGz+zxTTrgOu0Jw/AuMYgb+2MSeOYtozyNIDZT46mUzYvyPuwT
wNjp1g0nSMyYYY09K/uBdl6t5q3bKhIE+7YkCc67jRwmXOr63U2lTcMGiCynIOP53DqZu4PbAd+a
NyfR5B6oaTo9HKDocNYi5Nf+zdd6uzN29HRDONCy3GkDRqo3fAOUuPclwiODF0FGw1Ujp5dZgHgL
93nmWzyxTghF+YW4jYIZ6DKeKzbmFNifM9i5pjSoDlwRa6dz7j28mvseczuwFlALErn4tDRlhU40
tOCAUeuXXfYWYnGIqRoR83CVHrmoa8HngtmbOLYXdAnnwcR7X37IEhdo8t9AQgTE8H8SwYnoHE7F
Jb8J0JH7dFZrl74yJxI0msh3/MXIWzOwY9YmLymKoyRk+oySR+/g+u6Z7APk08x5nBFYrERidrfJ
pM6jEhCCVUvJenN8gv06uqeJRi+tgQDXVQAoChBMYk4ToR/Yp23HRV9BM2RB8QpA3kEtp8y7KbRB
i2Lw2waQK07tf/w2SKiKpBml0GICXPsxU4iQ9xq8hJJUf5neDz4Ai8PKmFhqCtC22MGHj6mhsWVf
wBRq0lpKkZo/zZt4s5yLQdIqAwHawDOFD/yaohj/SGfEWxoDYfbU8X5JbK/zyNVkn/2BDQEQ3uz0
ItiFiEmHO5t+okGNs1wfgzF0qUEF5GXh28WmIzWIal22fYaQLZGuBrC+lrLqLaKQGjH899oWNMAE
jF29+nFGHrGzSjEOnNer+EX1FoC24NLLSohv9Ene7Nfshv1coe+sFvdlUIEnyfvx01K0xTKS+6al
+eQMCU8iI5O25IdUXylNF/XxM4w3EPv68DLY0woWaUH4TNAcDx44rW8Znxxv8WvF/PdUxUWlY8oL
bO3jLiMelXEyS9QBi6r/JFwlsSEmuFFs6qPDQ+cyjX7S4Cu84qkovzb9tJO1uwWy9BQf4C7iuhJ0
+YyM7i74yFtCFis3LIvJ326+vaykAWRgCY7w3BvbWOsDDxMXs5r4FFDMO1dIYlgJv9taLc8nQmCY
0h5pawTuf//zBFe+3XkJSKI59DX2rOpNNmTKwH6lu7C3YEJOBzay4Qp0r38ZZgR9WF2B2/VXgOe9
/3IdyuNd5t6o9oevDa64nQ0cY592LPrvnewK0OcYyx9sK5RBxoTO+iIejDLHCnObr0uz8spEWg5u
eXhaeXXiCxCaLQ2s2nWRk8Vow79A2Ooe51gOZ8KQ3FL054KaQoV9XKtPnL5mADWUSiF9EiZPxl7d
aE9xlxWylxqkTn3t/ygQE6IhJwMryu5oheDxWuU+xyk5515gwbFsPDBNO9rZuzXfwr4khNfOr+wo
IyJMNRL5r1NlmDH04aLjhqLw0LsJnF+Tykvog+Uo2EHkBI97xb3nZU65JT0SpbldaEfcdFDyk/vK
pohZdwFM
`protect end_protected

