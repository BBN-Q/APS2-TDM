

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ncUawuo3vR1ZycZF8xtqqfVI6gCrdI+PWd72xdzgvbKVjiUqedCWSUEBFuuQDLCwTlT4hYrqtcoA
k+jkF6hUqA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
N3KVU8m7dp9m/o5klJahn6JrAp4dPvJ5px8Qjfdd/9teg+MgeqRSyR4a+nedbYovR1iG1M+OV4GZ
eedyUHeQwlftb33WHTgiSQcQOeDYQHOhB1q+SjuhN26SLFWK3YFERu3kL1tM5w3W0nuFqj+bXHZu
R4gQdtVWH/+OjyCytQw=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ZuxsHcVs7eB3t+mMECRU+c4tWaV00xKC1y8JMSw6ZK4lGIrGd9iKbAKZ3Blwh1vsVCQb3NTC7N3r
Y605Rnu1VKPlFpM556/vIzoPVRgcSvlo0qBj3oTSzlA5eJk5FVF3mP4v0RD6iY8xceU38ESPNbz9
tslYUbhOJVSsY7yCjCM7p+456bByCG6ed5+0nGONoXPAT0zF3Hxdnq8qgQDMjEIvOsaFSADZUSxL
WwjD6WPmcry72t5+zgCtiIUOoGhbFWqTndKP66O5YJAWE6dVlP4zMLQZZAfmdfQyazOsgs1uciSH
+eAOcN/r5BkNmFBVWZOF8biq4mt3PmniNwcfbg==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ygy9fvZbqToh8lhxP+oGEoqQi72mLbOonZqXDBQOfdz3oQWE3Hi1Zc2hfB1uR17TPoqAq2eJIm6k
q8c0om7asQ06vgODSHayDyQ+hyxq53TnIlLVx1AtJPfm0kI21kep00Mfc/Dwi7Qyt/ia2tlS/tQw
4OktcMlj77AyGCR8zdc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
mcqNli4YixoMqmYwzxOZ0byTQYAQvCZuCaZ7iJ4keY79GxqKVx5edvY5HqwqCRXfHCDzwy4qGKcN
pXmE+CGNG2mMTGEfU6W2QQ+HDW5dsb4d7quBuFh6+SnA7XZEst6UjKRr26YyBGTL5qgiRLyYbkFW
QKRK7TmdgdCAj37TPbTPR6zjrQ3PTlWUwzVToIPxndDd6Jgk0ZyBHqXveC/6PEihQuzGKgS5GKHX
85sYZQakcEpa7RtFdztUyxh1/Do/cjYhmERWgZJD9wSCPweFJCsvo6MP2JripEEkasaBYRqfxMPN
DPHGfcHemBvMggmA1I4jVeD0GpW65Lo9IxE2YQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4768)
`protect data_block
0uCsY2XuodQaeegpPLr8Jmjnaz8uMgEb2UJ21dCjokinwBKHUgbC/51IZlzHgRjjI/UzZ2xG1Rzz
OhqrrsHBW5JCsiHqCJsNKD2cIEzKiM9SmXIxfZ8JxhKNWlm4ELgiychgf5w8MTTUya4NNlOMeEg8
Zx0oDFE3oNCWwwxX10IbVmmRCIOO7vDBAjgr7l7P6w6PbGSFOlji1TUDE1m21RC9LMAdIHARFvJu
zn5v5eqNTfD1t6tFNZG6yoh7hy70eM8RhSjfsHQAuflERoV4Z2DMiXKu783uJ2pyvuNReXbGooiW
WmPJg96vwys07+MRAd1YZqNzHgXGDZmuZYtgv+iPsoYF0AdokOnFmPfo6kUJOwQuUJuUuqJ3m+FR
MyqGqyV4Sx4ZxIhuM2fbLWqiy1PYPkH1ns5kHDcm9nZqfrByJv2DeA7UF7nILQfxmdp1vhYfMneQ
RrFeNoWKun06RON4OikAW9AuVsoEbrgcyuw+s1gzT/2oUGDdZr14J0Z+OC9qsV/W7Zt9C0fxr7FA
CTUyzDSxhpvMJBTu6NCs2tcZmtYxWK0j3x9ZMV2AUr7zkAeCqBC13ZZmwf5wxXKldV5AiX3P11wy
idclLJywPulsu0lMIMN0/exT2uhTeU9PYxPJDLWIN4dN1OfdJSthAjPCFfRBktv4l6v7hu8VMAQB
28lynGijbjYXZpFZU1IWbc5W83ZOLDV9SuRMtTqU2aUlAaNY0MJ5+hBfrSgQkmDA98jERizzgIFw
Ppfedpx/v4rr5MzDvk5qamEtpnHv2degYYYoaG/C+fVjpdhG8E8qTR9lWMTxPkS4MyqJHEqFX/wy
YD8ZebKsMd9xk1ZLOJFURYHFr/M9g43BlsqZbjkUVB1JJYHE8u5LFxqmTVasD65YXyxPAHfA85dT
XyKlzLZ6x6XjSCs2MqX6722yV2tFIF2Kb2G9DjvU0HcVngAhe95lcfFZ2JWX1n0XVotS9QL0dJFI
uTtsk6luRvdWEvBgP8ehrcbxrzwLnO7QxXvlxTEFhjXXw3d28jSjjMZCXmyjFebiLKteNii/KNtX
60fCc7nZVfmrtY85Tjxjyij/Sis6vc1qZZBhZxmeIaFFw0ZLbPG3lGGd5bMgHCjQ9qi2hFE29b3S
6K2c2dE1dW+JoSdm9xhjiQvZGWNdKpFbF3iDJGJL09nQX1MMbC1iP7FhdTUb6HV1v1AsIXszjbUe
KnMmg1xyuACBxcnOAl3O7m5RBC0SfdZ7BcnKJZG0hg9wf7TnU+asuznSh/ozHbllQWBqtyUhA0tL
5nf6ngeoF3n0f7fUUq5qwkmU7J+QaBvcSlnuh+fEdyWpZwPHY4mEn52SmhvtVENmuTkiY/afFgll
99vwz2T2rB4ZuIuWAX9yRFqDz8/zlPIwr8er0S9tQpbmtGMs7U/uVBKQf6zswwMerhnjh+dnfAc+
8Zf7OYQ/BF85RxUXfQsx92Q+B7InaNWch5yKnR3KU6jGcGYQNfir/hN8wj8UHtml7Sp0q+QVoBiL
boUFZ/BMuXWEI3J9UzsZhRqi0TW+dqDxDF+csRkyD2E1inaJi7w1wuu9/nSgMTqqT0shFoGKiXTn
aTx6FZ0HBLKuBsl2UR7LW1H4bTjvMZmRaUOAfOrmv59bIkDNP5YY7zb6EcCZYMr4nw/PGw2YLDFo
j4z34MqnPn/I5KSG3KGlyPyoudjkfZmHFdF4q/I4SFBbSAfAy/+1/RD33joawjWtN55BKTluPzMn
4Oa5W6rGT9xIIDJXpCNQnBNZrVT4KxbtwVB96R2gwVDj7bddYTMoZ0IrnscCUivDLpXh446Guh8V
JBTYH1hgabc2EtKIh5ZcpJF1s3hN5R52L57vsdjRYTx/Bw779mZ2yeniW5FcgQSeDSMEJPDKEEp5
oHJ+d8MYk6Vp4ukVQ67bMV3Qq7NZMJJ2ZksiwWAdWf2PhiDnDV8RncKY0uyswIv+XJAIvJAhaYAM
MOstdBoQHU9li82N4MlqYaV53ppldZMpY8gndbeHM0Ncl1zl60vgR2nzw/aST6aJbmwYKpYMYalm
6+3IY+djBaELZytQI1n/Nnc2pkeDE9Mi9t2Uzh/dJdbV5BLaX4mX3wjG+pelAfjXaPLijaimI74V
JL8WihGVz5GRp6Yk8anRYkGKThHYFdj5Rcvw3mgfQpe/6FSYtDFi41f+77W0TrrICw5D+2YBsUYZ
nMivqsGeA853vqT788e2v5NXiWOlucnriunHR6eIZHKRQVx7YaPqPbB1e0olZ7vrbgaoISH5fil1
8qMwLveadUuTdo/tohzVLimIRnJnGKkjPQFkT5gl9JyB1PMisdlwSSdsWkuEL+EDuSyp+e0abjVQ
sHGf7bCgstquQE4Z1gZEW0XsVwNloWLwlst6IZvB6tuylJdp4irFymGOCqekoQKBJh7TP8NyLyZv
yMmSkJKZdlrO/36qORb3M217wRsSKZh3MZrnVRvNN7q8yk7QuRHrblvZv2YBnm//iWySMBr6JKEp
RZGq0NZhdSwjS1ivcDXjj49uG9RUCAanLwySQRpl1x4cn/wa179VgcyG6ELSeEE/YyjSXFhIlhBG
x9eUvDysuAhkgfU1x17UuOKuc/GEtSLtHPDcidGaWdYySHSKRb/dtqfJL6CZI9YeN6/G56xtefXy
6Leyqq3g78Nh53z2Y6YFlfsBdjO5oh/9sDb0LvCDWoQh+Ll9EYUwBolkyCTKhc0UVNpUvlZag9O5
w9aCN7wBWsMUsOePfALWBm5LMK+t3bWI+78h6aH9gWHW/pl2QmD+cd7PMsFV6KCRbGM+SiSTwze6
kPum36kG+CabNKqZTxQ/9zCW5YsW825VY9ZYBeIYcqEsX3RscHAnyhskbbZJF5G7RRik9OvHY1kH
eGXWG/ybRNMAtEnYIm4R6HaVUO4ztrLwvu3NtBs1jJFyg4n8fENMahY2BZFFsN7sXXYweGw+/oNl
T4/ZuBnPc+TtiaalZ/5GNBhMRkARLuE1UHUSw5TM5CnoYnakH9tplHile2YUFcjtZoCEJ5BOX2Rq
V3D8YLPwaajXS1anOXyo0zv/oySC68NapkhCAG0vVb2mjB8ALLW2ao2ZCGHcx+A1nxnAhHsrtjhm
TlYXxCjPQ7YXm5hWT8Nkcs+MfbT76BQMYxzfFS0i2G0Ih3YoclOgxutAJhI6bxakX5kojBDeNto0
rRYMVcvYAgD9+QYqPSPT3JAEUtkzOzlGN4UjsO+u9aFhkgKHiYAfL2b7MPrNKQ1rNhlihSJs/0L6
aGx4WxGknn+6qVt60RRjYgfHklTMhtuC4Nc7x6Ye3KXL5u3tEhSLzExhoGICyna9xoRKabyIAp5J
sJXuQgDS+DwkeDJ4U6joG59Ow8hbqBQLJRzNvWNGv2df3FBbo5PqxU6g+1k29JXtChuj1bFQi92J
kjUeOiWD5OT9NEXKD4mIKLBq/XQCIcYVY9ubWT89012o2jD4vB6VbSDwu8xIG/bvbLDvpVro6DLm
hx6wBVNaPVgIo8gENzvw1qy/5bKcIip3TLWOmAiv06JLjkV4h6GdhvqD5g5m1M/tg4/D///Ir2bM
nmvzInK7Zz2wK3S/KPrUSLbXikPLl7JUJuB78rF6papjeV4Kau8b1yS5gPpbKg0D1W+7Y4aSFFk4
g0fZQZs7+XaCyibWrvKnqZZ8Z6KqgjDdJgrO2ZA+7ggEVsZIwJq2w2QXC6UhtNDNGPHuh+zS5byr
LyCUZMkGDoAPwCX65bK7JMayADeHn0gV01X9jfpFIRq+oKETtAfGJgLtm2OD60ttXNRCTVzuoSsS
V7B1uZzN4C7eImrS87Xc9+WI9pqYeOXijsrHtjwmlVRITbMQE+m827EZFwylj0WrjF48kqTlNFeS
d3LF53sdUUomdKm+It0X5hrPH016nW9GyfRU8ZlaGnXNoicKHd9I3oouFk0Y/ZdtcV4cFqu1I2m9
VLm0mSyhOKSJlpm8jXELMtgvS4AMvL/opRJu21/k6nfi9PJzLgqFhQc3Y0x7kQoyEY6WZU8lnCZr
TrT+dY/g8egpko1POMK4k3cvZyU24UfyFqfdfLQT2WW76m0kEYQJns++u4wXnFXAXpy09hhas7EI
NF8V1xUu5Kwd7ZC8Wvosj/gU4wgV2BLLG4Fp/SEySALM0NDN9HjKxE7ilELw8kUTPgmw6Cr0Fzdr
Dhx8fs3jOqAi9W6ICEeL/a8N/vIKC8OrCjgpCbu/bEME4bQSrwB0lee8q5E6QkncPM/K4RcB0L33
RdD38hBFRoP8YiZ56NocECmz50EnjDFkrCEUZIh9SqXBgL0GrDBYKzHWGqEmfFWLzimXr/G82YPX
TL9tb+LiqetCUCTEW0P2Wflp73DLArfMjJ8KLDL4ATUGCAMTbHScE7C4SMq4XFlMEeO6O74gDwB+
6YSBpd9zFQsYZ6XOJYDR/U42Xv4rXWjG4HgmiYWawaGpJbIy9YI6LvVX7aH3AdQ5sTgF/8lupTlD
ZwXTCEVd3768SXrzYQfsA8AJADFgJHWeBpFzy0aPUpiAqnr8sq5/Gsc1PyD3AMfHqrjdsC/0HQwM
uHSvqwyJNSz2SKgXia2049f44RH/2NApfFFuJsdUewgYmM0DwyG+wADVCvrxhU8k8ISPvc8kseYF
lI2DqHJX0eL2G383t/xeAADVLvH5pqqtjdVu8icVLFax1A7lGbPsxybazGyy3/jDFcW43zYJFXZz
SvQP6JBqEKel516UpoDAtaX9pC1KBHP3EEZaRWCKIE0L95VaY9aHgeoXL14lY3kIPh+FPDeBvLc4
QXUsr6bmzi0GRCOtVf99LzKERUxpKHj0foCcLwpoGeIonn/Xvg0/PvhRaVcPnE6lA7ZFWn+jsnW5
bOmSUG+n77Y51zippf5OSpopdPXHnMW0p4qXcQOpZtaDbDWhHemgopDIHF6dY9jsvC8ifDEpIwYV
yJjyN+6VribGqnZfdRz2Uee+yRJUjxb9j/fKCTi/y8yQOS9HFTVlWEn48YbJfnKRJwSn3mmaDegt
04zDI9PippHNXGoSgiXCQPG9X76m2XjF8Oe8pGoWz7Wf0IC6vUiv5yJfbZ5KozHA/DgU1Zwl10tj
bG561bF1ZSRysg0NOlXXeVfHYcPcyigljWcNlMuZ2hjaaOTNPt9BvnjHAALjYDOTwU8B6BRp47vh
UygzaTvaj+e/LnjaeKpsE/n6C5KI/bQKHJjjn/e3RvXFqc8YqPi2NaUctW/ebaluQWtaJcCh7oiL
K9DLRYNrXfLze8S2e/CYjjgBLGAHwhs9W3S+MUUtUmUWrBU02KXmQpdCgR2CnF0wIybXd5djOfyx
sStUZvX/mpdAzhwcm8t4gSK0Yq+kIY/1ihjTHNrbdiCqXBwS9747ZkQ08CI933ZaXKQPGJJPBvdp
bvSbGPgptQVvxg6JRD3cYT3v36KuC8GItiJQi7YKsP18oqUg0P0INty6aTjVOmFN6u4Ovk6WCj6d
ELvyQRCvyNlyW5/IwbJMZkOuPf/+0TPvuZbnRRKZUP1y0qK/Xrib42ll/y2fPh+hqp/LP+YdTI/v
KeIn31IF19i4w8uHQB4IwqVSjW7pfYBTqlNIJfbBssInZNGT2oR7FIYWTiFM7+/JbycF2bzM5u4u
EySQ8qCgoeKndoBosqb1jacdbhTbuTJTnF6699Os59pqjo4RHuYvRW4455zfoC+wxCrrsnoFcfwn
SXrfIi1fuxf9oufL/iSUJL06irYpOjZY8GtPrl/MpgQLsTN0uaK9LU8bJCrTaDuaofGsc1ze4Cgy
jHCsJUvVsyoBzvP0jXjp2DVYw5yDoPX/Xk+2xHpCCKBYlzGymkG+z1c/hE/8n0b3SYiCQ9joOZIv
+CaQ9wVMozs/dW+J/JPZmpa3dMgRV0VAVnYyJWezm/kUiQDForj4u1TcRwyTFOM8cG6nmhGezsRC
bbrl2AGeIAiRYgJlxfOW1XCs6+sFMv696bUyMh2Q/WiIW8QRMSmsjL8z9brmqrP9whZ1rcjQFYN2
VYEwUeXrk0uT3e+87GIjn2DJvuW8HZocKRroo6jFekgYi3dkYWewONHuHhuGQO6C7CYtzlQ2HKmr
Eu9mYG3l59V4VfFt5MS+VLEjtG07YrcC8/65OQPD4B6YkKZrvDH//k1jQbGlyCSSo6tb7a6ZPBbx
9/mu9472dmpu8KkBAjtmFYtTEU02GcbBQ5HYUl4ZhM7gas1j+ZZGx2KfdtQD0LTL6RdQUMmIhDUN
BOvZulchVSPaA06i1S1APL3ZrU4XNme6Qn9r/qHvXogub5dnQvTEtqITk/2pJkSEsYLbD665DOYv
eVEc/vdlcljsWfDAkomtBft+GN05lsqa1nAMyEeqcoX1S2E41w==
`protect end_protected

