

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hIBbF+kq3oVaBXwt2/thZmZVCkqEUsrobKuL7n/Is+v4/IAZD+ZxnU18s3JR+GBgEFSO05ZDR/P/
xVqnh5V4xw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
mFrbrNN2Iy2aMgLbmjyLagVGv1BRA/A/dAXtgEZvBXH1JsdW0tbqE7CcgD/B2t/bWf/vphzdyEfE
Qtz1a+CCHs4ZBStfoFAa0Kk2/N4AElHqndo2m2qkwB10dpRxHYBYIM8TsnGzjHv+Gc3MRRv5nDTU
c0fluXo+oor8ssR25QE=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
DijfY6YIFcLzBTBsFWeeH4jYfY8NXvmEK/hZQ9aT0hDSd3Je/Yj21LmilPHhv70y1trouG4tZlkQ
XpgM4Go6KW0FBpBt0/S2a5XkCoVlqKCnoc//o4WuX1mp91+H+1sSGdHdOtSMW4j5N7yi8fdf3Mma
iaJg/1V/iPoZ7fsaYSHM1whghXW3BgAg+uVNwDgKp0Xvr0+v0TXEnhMcvfJGCk7ZxZWk2u7a5iEO
OrSkH1tRBHn9Qs31Uoph/IE2TzjfOAWzb9vhqVCkYjlawx+iuHQsXxJdeZzjNlXERo16SR5o2JLI
GgcU9rsEUp+Hcxd2JjfSbszpWRHEU/3MaVNDkA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
XNCwdX+l36YznBeQn7kiJlUVYGKrBB2zjt1UpGWFaIdIOQWhZL6zxzyLVbRsejTTuYPFOE64n48E
kMQtjnzPGZyr2W3R3SGB6KeHHUx9pNxyeNUyrOXfxd3APJdAnl9DigbPc/K+n0zkIbqWEydLVfIg
khTPlA/ncexRV1pXoq4=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
P4vVw8BLyUspYO28urZnMeeAl1C8jySXctEPFVvNqtg6Ihava9NSbOfscJ+47pmoPKhiyUWcqNJe
xZD0jdlH7PDpmGu9W5rxevvgidGt7SMfg0iUPqEmLLxZG6dlkSkZQKHeBdCxVW1l5LVS2iogdVV9
APcLIH1Hv8ySZWwT7HFfcdud0XUs4SZwhceaZ8TiRT3yp086kneb0uW/2QIlfzI1uwVMn4U5QPIP
rt59lNQNLmXYEhGyXeiqJ4sjMbP+3IG4yIeOFeDMhWUf6qgDysc+rBTvTouOsEPHvQarXNA7RtYJ
afWxcLBokJDKrgHjACFrQmNY1MmJtQUikTUFnA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4016)
`protect data_block
PY/uOioAAAABAAAAAAAAAPFMxADosNXzqaU6ZZ5rzDCnxaW37Ad3acEY0IIchL9MPE9YibAhzvXy
aqLf9PjkFWm/tQbyDy+YAVIO+g/0ycysOhYmpPVoNh75BIlyCUbafwgGYiHzkhISq5grPIojoXIB
yGecR3YAp+SVZB9kwnIEdG3DBSJc16FqYpHY9cpy6pjbjSzF2I8NPSPKzG+30s049puSRiAYdRW+
plDy4H0P/TqjECuyeJlt+QjGmC3uieG10nvO3nNGlOaYCFjRqOiRmn7pNSnGvGptqwFY4jh5i8Ux
EOu49y2SUFcU3fX0GMrHpsyGggMhBKcX1m20iSjSLdj46JThj+ikP40o07nS6Fm8sDUojO0K/qDa
HQtVLRJOvEpRpOd+AwWHH8kQtstP5dQK4UlQUB7/HEUiiqQlNu3yL1zKB31u9A4O+V/IsalQ95xP
7ryxI/P4kwHybjQ/zRUTYxJQIG2pQBo3QIMdQm0EmVu6F+sd4S1pqMlUL7yblwpKlrHVnpwj62cy
uy+rK25cokyyQ1cVfeQR5VH1XNSz9DEnYHH6fQScCYX4Gfml0wGjV0GgYyPOy/KgvvGcbbfJBAi8
xPv7ppQaipkBnHIVzrrFmzuL9D8A8/rvNeXep6wRu/L3RSDw7R7mIYAueIo0GNWOg2RJ2b3UKZNV
c4mzC/UAEGcZi8cRf5yy4DqC6MJoMWJGhroUkzUiCC2o+WTnpZfq5eEXKqR6e6rllf7zjrvV5RjG
L+o1fzG3m6Qt/Oaa8/lPHTSP/eqN7Ma3YbXIuWVSQvgtz55L4qE308iXTzsOuIRnwGP5N7hLL8Vz
ZuwnNwjwk+xKkj6qSdwlq8V3kF6RAj9VZezy+Un8v4DWP1p+0WXVWK0WsZVWTuGBxB4F62mT0Vbx
xyz87SHngWwohTNKW2gamfxdYVNq9cCkI3/hSNDbumfFeiML9lq78F9huiH059s+sfF4plmzux8I
LvcCWaZ/Jve+LhZcyVsGPNt8tWIqDtOH5jkWSLFU6ae/e7NcizmoS3eerbeZwQTAD0VAmDD4Iy4k
zUJF0VwNj/vx5qJPvZ8sxbWuH2R9UE1SRbIXJ8hKYgGlzVc0hGj3MTUoCBYhc7gqD1m1JideMx+f
AJZgAv+yb22VZ0BdkiKL8JCz4wo2dbMXVivoKsl6/S/eu5JICeUgV2u3uhGShWNmQQUGdCAocwYR
vRE4KhCCyYpgNwW1moGOUZGy1WZFZXQ/odrsS4md30riW/mu+d5w/gCYj1N9GywZH6eG4kiWRrN3
lixQp0pdxjBTS4m3bfj3tL7HtGMZpklxRSVvzrVH8JH05h4Hu7a/4bykm2NkyOZWPYBGrgiClliM
7lwobd+xz18rWu2vmZUodwstzyhV6wVopRd//JBFPk4x+br8VT1dpOBGRGbOzallEETIPmOG5pa7
mrB8dUJ7Ye3tNuWK570VXy2ov9RYSwgA28Psh+ae4dKeQJ3E9N4jxwxlvO8FSt0dG2gQEpyRVnRH
hAFVbkARNTcBD07oiuS1YhdzIFBfmdLY+bGq0aWR8O8jONW7sWFW2q+WtthMgJGcXE4QgzICgLFl
n7vUHDg7/WzrgeThzboKs/MPMMZ5d80jtihzEebZq/WXjN01wNF7ekAKwq4JhFuXfMKaSNF5aMoa
tueowQWhtUa5LiIBN4GuBpFKyXmdx3zY9VZMCNKjpEI2TEgfIFFw7kqFhajyNji0Py7rRQlCJkSv
oKk8rVhAIKcMcsYgfGxOIEDBW0Vc3l4EzzY8RbO9SERNfb8FRbsWpZ2TO94DRZ218AzWv0J0FUtk
IlmAaz4u5UJNt9p4p5ILjiKXcuIcGNGmPx3KW4UiRp0xZ3Dbn1LXQDHO7eykUxMNrp/mRMAFI8iR
IYqvZmN/vr81K0QOvnV9q56K6GtIX4nBumxReePiBkx8G833MpTyPRp+GMzRR+bBYCQtplBr+/bD
5PT5cE0F4q9gPti+qXdr6lNghpy+uSLffxYFxMxyHFiRg9XS1t6GIvd7YfocbWFLZ1kogq13MrA5
kclNTE7E36e82QrJBmJX/m39fVOVy7fkF6WQufwvFwTPlj91sMcTiWmC/58Jrd8Cwn+VggtTCXfe
obs8x4rLfbsfDSUmy5vU63qDYxUOhwGhZOkh3Wmodep8gdY4CvKSn5Ia8MZvkWib5k5JeAPnuY19
rHsEnq7DPUtEseUEHboOOYxWHkxXdpQKc2ue9SvOdHeCo51jEYs42BMVwpxOLpB8hbbhPxYxsZpT
xAr1mN2RrzBtLp+6BlIwU6XkgDbkjg673Gk0zzSpY97tBvIkpVBygOFHMQ/yAPC5jRNNv2H0y2KB
A+l6AVgA5317Awr1fUkhk9JEVKFJxs1Q0bh7yYMS454rmGxHEalVq1Exq5ul+GHL0H78Arz9lowj
7T+ut25UREoumY4FhlqCzzkmln2pjIu9+2CpJ8I0YqwezGx1aj0vGQl9eHRMy0yAS3rG/RqdeFB/
ybnIk9ZQDxztpqHka0cfApQrPo5r/LA6cFUiG/6snFnidU6KowzdMU99iEIcHVVa3k1KoJHNYEue
NnatvIiIC7sZIci57nKqBAlIjNAIynT5XJlcv/dITQvtPbH4HVxM9DLTwiTWmGz1NS9wKF7krJrj
xSOC7/JhyiCS93NSFLLyzYZYvaFkfS26rfFAbItd6JmKAXdawI+m59Rx88jBo6jKNGmovlouoltM
ysKZOiUsHZyapoDdeIf+TfXRgJsv8X/XeYFflY2lm798hmtkh64uAafjJfViPvo7+cpxGAxRuqki
GdVIweRuT86lQK/DmELQ/R/8sz0e2KIQEoydTiroaixtJAa/FEnsLFtuplyUQbS0zbx7LHwT1Y1q
XajbmdOlYhrgaevF2sZm08ev1CNKd39TDAQ5+ziK1CaJzrT7BJmaJV/a48vRmcpWevipSto6Zdjq
O+eLb8+0DUbFS1H+tD4AwlLZO1/IpWVoaYqL40X9al4c2EXnEmbnWgSy4o0pEGaAumt64rl7J3Qy
SKVotlsKYejgUjBVLfVFfpaLP1qPTwkdckyutjUDf+begWTlYQdch12946+X27c9E8LHTM1iBPCe
d9JXZQA3mQ4woocrslFTvuhmr4DCGQK/MIJkfZY85Md+bwhOK4K5Z3LqbvTBs5EzEg7m840b4cII
i3eetl1rGgxj8+t4X/NWrn2u/3jdWrmQJWLbkQJZ0zVPwhB7CTuahNQjLL1JjIppE80JOrAo22j+
DsbLVCjCIwmycdTWgIKkaDtQ5lP9gqeDxkNvx/EItcPkNT79E4dSRGvWVapUCq5PYoeldr04J14z
ifD68J9jz9hDbiQX+jLlBdt04i3LNc3HMWFBlH8QdDDf/gPY21lTx+jaiOPqeMhO+NExm6H2YlPj
emjjkznfyq/EGPD2jfv4cQGqTJ7WOG5RlDUjOnit/t9/XL6MPXPgiSQGebWP+lFHO1NwENZmGywO
+Knpb7OPsYoZj5WpTIK1HTjND5ovUQ9eYXpMKWQvYF4qB9ApNezxrleu0WWeCCtmyy6MYKjZb4lI
gWGsZGCwp8DR/jVS9rf0rWpzzt4H5Qcj3UNuEoa0CS3ztnk821YwkvZ9cOEvd8V+rl5DfnqrqiMA
1peBt+gYMd2Jz1MrCR0nsideRf6Re30+sXq3Mq0Kji4RumFU4UUbQ5C/2O3B8tvTGKcfRTT2SBg4
AbViL2EL4gY9ut565OLkpA0srwQTwMFfhAkMp6fsE7BtmzTicRcu+ADnheiujJPgePPSQz6Hk0Do
aaVW3dSuORUNT9g5/eViAcLLO/QnZ6/r0hFttR+n8VGgHOQaYCBF3NV/cNpcJXsk7+kw0Lu6r/mF
wNrohlcDDhzTN/+ULVoIvLPh3f1v+gxi/Y9pwD8SYsrPQ43ubNYwztuCS51F5tYPPZNAu+kg1xLO
iV24EJyYnoKXVWFS/pypWnDtc8PJQuOXEogDJDsWtqRyshZaDI+NiLwq7AK48C/o1AYA8Zr7Yqsr
MlH335VRMYyNdIOvtUAqW/h819Y5BTOob98mTg1fT7Utdw46xsoXNW17cws8/TCAM+3GnTTu8OUi
uQbRpLen6vJHa5lr2+zpCVQpsTZNNk0eqjJnitsMWoIBi1ZNa7+V2LoO3j1WPDXqbV8lwKVgahmA
bfUk5LgwtmHAKunn716IeWpsJqtQ3QITtjfGsB7I9pOglD+aVK/xcOoNCckTGPY1ncqqehAIoqgk
olf4L2oS2WAaEyxOBG/QBVCb8C8U3RlZAPlZbeJ/aocN10XJnXywFZfcToIdDCWBc9pzdNvF9ujW
Gz6XGwwCV6a0p61vcdYMihUMj1HG5nlmQX6RlCa+Y+qQm/8cRlqwf/psIsk8B7k5qnJzXnW4KYwW
GVGgA3WMpMmwykEnJqmGJuesUKLDLi5VI0YxRCg1kXyP/KrpkzZXs8B4jTXaxqOElXNsha6B/VC8
5E2TtqtppnEkwEFCeOnRVcRP2WZr1JLnYONZ/pG6vfiKpS/2nDLkXW6GIVtR4MbLQOf5XXSeur6Y
5D0kAfYVWLXTd4DHc2I+Yhtr1y/v9QKOiwYlDi1Y+V9U0Uz8onInNH6If70CtBvXWnsqFujcvMyC
LEsaIEB9IPszs7XKx/E9nsaHu4TTQmRop7Uvo3p/cocN+rChYa30yvRl6cgLI4NuBa8u9bmjWUnt
he9Cl0sjcruVRwnb2JRdhmVHcK8h5pg1220O8tHaMiEKtz19wHYAQ4d4YZ5N7qhTlMflA7t/d5iC
yz67wvRjyXa1ZFyhLi73DXidiGZ/WqvjAQPkH411Cjgh+oou44BxJu2wHFuHl5uGk6HgUUAd52g3
Bspcb/YxaalbHXgb7jmcmT3TO7dLIFQul11WZNBgmvIExcbUJ2TXNk92ANaZ3O5vJD7i3Llpn2FN
nWsFz/coI0ZkN8YMMGCjttT+r1inqTP6cj0s68Rmtx5FOAQeQ4zZorL0V0uLQfp/2SU3R1D9PSNv
vZ8HpxBSl+b2V8b7OqI9m2c/GUNi1IvWoYPn+46r9w4vb7JmBlFg5uHbZgMqQ3Q9R+bDCJXygq10
RU0uCYBgWt5EB7ehCzRxdMDrS7xWIMsjvUiymkR3zq6KtUwjPPN+LrZYn6bBS9lbgS+/iJ2vY94/
2lTXmilGJGAdtQglMub52EQwfAEcimcrF851ZUzD3p0JkcGuFlQ024aXajUH2Np6bGv+fzntym+1
FfP0soxEFWj7nAgGl1HPG8BPx3rj5aEqYDf6I0NLsLwXtBZXoU4kXTUaIKNlmLLpnpn7pMkt0GOK
/gXTBe1qAIuiXtmGVdvgWMcuHWpWfw38vao=
`protect end_protected

